`include "para_def.v"
module stage23_tb ;
    reg                                            clk ;
    reg                                            rst_n ;
    reg  [ `MAX_ORIGINAL_DATA_BITS - 1 : 0 ]       d1 , d2 , d3 ;
    reg                                            m_en ;
    
    wire                                           message_en_out ;
    wire [ `packet_head_data_bits - 1 : 0 ]        packet_head_data_out ;
    wire [ `fast_length_bits - 1 : 0 ]             length_fast_1_out , length_fast_2_out , length_fast_3_out ;
    wire [ `fast_message_bits - 1 : 0 ]            message_fast_1_out , message_fast_2_out , message_fast_3_out ;
    wire [ `packet_ETX_data_bits - 1 : 0 ]         packet_ETX_data_out ;
    
    stage23_encode_module stage23_encode ( 
                                          .clk                  ( clk ), 
                                          .rst_n                ( rst_n ), 
                                          .original_data_1      ( d1 ), 
                                          .original_data_2      ( d2 ), 
                                          .original_data_3      ( d3 ), 
                                          .message_en_in        ( m_en ), 
                                          .message_en_out       ( message_en_out ), 
                                          .packet_head_data_out ( packet_head_data_out ), 
                                          .length_fast_1_out    ( length_fast_1_out ), 
                                          .length_fast_2_out    ( length_fast_2_out ), 
                                          .length_fast_3_out    ( length_fast_3_out ), 
                                          .message_fast_1_out   ( message_fast_1_out ), 
                                          .message_fast_2_out   ( message_fast_2_out ), 
                                          .message_fast_3_out   ( message_fast_3_out ), 
                                          .packet_ETX_data_out  ( packet_ETX_data_out )
                                          );
    
    
    initial
    begin
        rst_n = 0;
        clk = 0;
        m_en = 1;
        d1 = 264'b010000010100111001001110111111111111111111111111111111110000111100001111000011110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        d2 = 264'b010000010100111001010011010101010101010101010101010101010101010101010101010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        d3 = 264'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        
        # 100 rst_n = 1;
        # 20
        d2 = 264'b010000010100111001001110111111111111111111111111111111110000111100001111000011110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        d1 = 264'b010000010100111001010011010101010101010101010101010101010101010101010101010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        d3 = 264'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        

    end

    always #40 clk = ~clk;
endmodule