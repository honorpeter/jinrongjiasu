`include "para_def.v"
module stage234_tb ;
    reg                                            clk ;
    reg                                            rst_n ;
    reg  [ `MAX_ORIGINAL_DATA_BITS - 1 : 0 ]       d1 , d2 , d3 ;
    reg                                            m_en ;
    
    wire                                           message_en_out ;
    wire [ `MAX_MESSAGE_BITS - 1 : 0 ]             message_1_out , message_2_out , message_3_out ;
    wire [ `N_type_control_width - 1 : 0]          N_type_control_m1_out , N_type_control_m2_out , N_type_control_m3_out ;
    wire [ `message_mux_control_width - 1 : 0 ]    message_mux_control_m1_out , message_mux_control_m2_out , message_mux_control_m3_out ;
    
    stage234_module stage234_e ( 
                                            .clk                        ( clk ), 
                                            .rst_n                      ( rst_n ), 
                                            .original_data_1            ( d1 ), 
                                            .original_data_2            ( d2 ), 
                                            .original_data_3            ( d3 ), 
                                            .message_en_in              ( m_en ), 
                                            .message_en_out             ( message_en_out ),
                                            .message_1_out              ( message_1_out ), 
                                            .message_2_out              ( message_2_out ), 
                                            .message_3_out              ( message_3_out ), 
                                            .N_type_control_m1_out      ( N_type_control_m1_out ), 
                                            .N_type_control_m2_out      ( N_type_control_m2_out ), 
                                            .N_type_control_m3_out      ( N_type_control_m3_out ), 
                                            .message_mux_control_m1_out ( message_mux_control_m1_out ), 
                                            .message_mux_control_m2_out ( message_mux_control_m2_out ), 
                                            .message_mux_control_m3_out ( message_mux_control_m3_out )
                                            );
    initial
    begin
        rst_n = 0;
        clk = 0;
        m_en = 1;
        d1 = 264'b010000010100111001001110111111111111111111111111111111110000111100001111000011110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        d2 = 264'b010000010100111001010011010101010101010101010101010101010101010101010101010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        d3 = 264'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        
        # 100 rst_n = 1;
        # 20
        d2 = 264'b010000010100111001001110111111111111111111111111111111110000111100001111000011110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        d1 = 264'b010000010100111001010011010101010101010101010101010101010101010101010101010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        d3 = 264'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        

    end

    always #40 clk = ~clk;

endmodule
